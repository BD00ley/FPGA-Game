module VGA_d(
    input  [(8-1):0] DATA_IN, 
    output [(8-1):0] DATA_OUT, 
    input rdy);

//TODO: everything

endmodule