//top level
module top_level(
    //stuff
);
