//standard spi module
module spi(
    //stuff
);
