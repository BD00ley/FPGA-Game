//fifo for whatever (row of pixels idk)
module FIFO(
    //TODO: EVERYTHING
)