//bascially deals with external memory from AT25SF041B
module memory_controller(
    //stuff
);

SPI SPI (

);
